interface alu_if();
  logic [7:0]in0,in1;
  logic en;
  logic [2:0] sel;
  logic [15:0]out;
endinterface